interface aresetn_if
(
    input aclk
);
    logic aresetn;

endinterface