package test_pkg;

    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "../src/axi_lite_include.svh"

    `include "test_scoreboard.svh"
    `include "test_env.svh"
    
    `include "base_test.svh"
    `include "rand_data_test.svh"

endpackage