    `include "axi_lite_data.svh"
    
    `include "axi_lite_sequence_config.svh"
    `include "axi_lite_sequence.svh"
    `include "axi_lite_wr_sequence.svh"
    `include "axi_lite_rd_sequence.svh"
    
    `include "axi_lite_sequencer.svh"
    `include "axi_lite_driver.svh"
    `include "axi_lite_monitor.svh"

    `include "axi_lite_agent.svh"
